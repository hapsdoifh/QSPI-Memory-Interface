`default_nettype none
module internal_transceiver #(
    parameters
) (
    ports
);
    
endmodule
