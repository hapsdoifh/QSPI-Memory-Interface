`default_nettype none
module pmod_interface (
    
);
