module moduleName (

);
    
endmodule